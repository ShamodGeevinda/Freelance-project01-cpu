

// module read();

	
// 	reg [31:0] instr_mem [31:0]; 	// instruction array
    
   
//     integer i ;

        
//     initial
//     begin
        
//         $readmemb("output.mem", instr_mem);
//     end
    
   

//     initial
//     begin
    
       
//         for(i=0;i<32;i++)
//         $display (instr_mem[i]);  
        
        
//     end







    
    

// endmodule

module OrOperationExample;

  reg [31:0] result;

  initial begin
    result = 10'b0000100101 | 2'b10;
    $display("Result: %d", result);
  end

endmodule


{instr_mem[          0]}= 32'b00000000000000000000000000000000;
{instr_mem[          1]}= 32'b00000000000000000000000000100011;
{instr_mem[          2]}= 32'b00000000000000000000000000000010;
{instr_mem[          3]}= 32'b00000000000000000000000000100001;
{instr_mem[          4]}= 32'b00000000000000000000000000100111;
{instr_mem[          5]}= 32'b00000000000000000000000000001010;
{instr_mem[          6]}= 32'b00000000000000000000000000000000;
{instr_mem[          7]}= 32'b00000000000000000000000000000000;
{instr_mem[          8]}= 32'b00000000000000000000000000000000;
{instr_mem[          9]}= 32'b00000000000000000000000000000000;
{instr_mem[         10]}= 32'b00000000000000000000000000000000;
{instr_mem[         11]}= 32'b00000000000000000000000000000000;
{instr_mem[         12]}= 32'b00000000000000000000000000000000;
{instr_mem[         13]}= 32'b00000000000000000000000000000000;
{instr_mem[         14]}= 32'b00000000000000000000000000000000;
{instr_mem[         15]}= 32'b00000000000000000000000000000000;
{instr_mem[         16]}= 32'b00000000000000000000000000000000;
{instr_mem[         17]}= 32'b00000000000000000000000000000000;
{instr_mem[         18]}= 32'b00000000000000000000000000000000;
{instr_mem[         19]}= 32'b00000000000000000000000000000000;
{instr_mem[         20]}= 32'b00000000000000000000000000000000;
{instr_mem[         21]}= 32'b00000000000000000000000000000000;
{instr_mem[         22]}= 32'b00000000000000000000000000000000;
{instr_mem[         23]}= 32'b00000000000000000000000000000000;
{instr_mem[         24]}= 32'b00000000000000000000000000000000;
{instr_mem[         25]}= 32'b00000000000000000000000000000000;
{instr_mem[         26]}= 32'b00000000000000000000000000000000;
{instr_mem[         27]}= 32'b00000000000000000000000000000000;
{instr_mem[         28]}= 32'b00000000000000000000000000000000;
{instr_mem[         29]}= 32'b00000000000000000000000000000000;
{instr_mem[         30]}= 32'b00000000000000000000000000000000;
{instr_mem[         31]}= 32'b00000000000000000000000000000000;